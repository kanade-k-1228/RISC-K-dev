module RK16CPU (
    ports
);
    
endmodule